** Profile: "SCHEMATIC1-Proiect1_OpreaCosmin_N18"  [ d:\proiect1bun\proiect1_opreacosmin_n18-pspicefiles\schematic1\proiect1_opreacosmin_n18.sim ] 

** Creating circuit file "Proiect1_OpreaCosmin_N18.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../modele_a1_lib/1n4148.lib" 
.LIB "../../../modele_a1_lib/bc807-25.lib" 
.LIB "../../../modele_a1_lib/bc817-25.lib" 
.LIB "../../../modele_a1_lib/bc846b.lib" 
.LIB "../../../modele_a1_lib/bc856b.lib" 
.LIB "../../../modele_a1_lib/bzx84c2v7.lib" 
.LIB "../../../modele_a1_lib/bzx84c5v1.lib" 
.LIB "../../../modele_a1_lib/bzx84c5v6.lib" 
.LIB "../../../modele_a1_lib/bzx84c6v2.lib" 
.LIB "../../../modele_a1_lib/bzx84c6v8.lib" 
.LIB "../../../modele_a1_lib/bzx84c8v2.lib" 
.LIB "../../../modele_a1_lib/bzx84c10.lib" 
.LIB "../../../modele_a1_lib/irfr120npbf.lib" 
.LIB "../../../modele_a1_lib/mjd31cg.lib" 
.LIB "../../../modele_a1_lib/mjd32cg.lib" 
.LIB "../../../modele_a1_lib/mmbfj177lt1g.lib" 
.LIB "../../../modele_a1_lib/mmbfj309lt1g.lib" 
* From [PSPICE NETLIST] section of C:\Users\Cosmin\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 14ms 0 1u 
.TEMP  0 25 50 70 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
